`define	MUL_IN_WD	32
`define	MUL_OUT_WD	64
`define	TEST_NUM	1000
